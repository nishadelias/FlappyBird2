`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:30:38 03/19/2013 
// Design Name: 
// Module Name:    vga640x480 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module vga640x480(
    input wire flap,
	input wire dclk,			//pixel clock: 25MHz
	input wire clr,			//asynchronous reset
	input wire pause,
	input wire [9:0] y,
	output wire hsync,		//horizontal sync out
	output wire vsync,		//vertical sync out
	output reg [2:0] red,	//red vga output
	output reg [2:0] green, //green vga output
	output reg [2:0] blue,	//blue vga output
	output reg gamestate
	);

// video structure constants
parameter hpixels = 800;// horizontal pixels per line
parameter vlines = 521; // vertical lines per frame
parameter hpulse = 96; 	// hsync pulse length
parameter vpulse = 2; 	// vsync pulse length
parameter hbp = 144; 	// end of horizontal back porch
parameter hfp = 784; 	// beginning of horizontal front porch
parameter vbp = 31; 		// end of vertical back porch
parameter vfp = 511; 	// beginning of vertical front porch
// active horizontal video is therefore: 784 - 144 = 640
// active vertical video is therefore: 511 - 31 = 480
parameter bird_x = 240;

// registers for storing the horizontal & vertical counters
reg [9:0] hc;
reg [9:0] vc;
reg [9:0] bird_y;
reg [20:0] counter;
reg [5:0] velocity;

initial begin
    bird_y = 10'd240;
    counter = 0;
    gamestate = 0;
    velocity = -10;
end

// Horizontal & vertical counters --
// this is how we keep track of where we are on the screen.
// ------------------------
// Sequential "always block", which is a block that is
// only triggered on signal transitions or "edges".
// posedge = rising edge  &  negedge = falling edge
// Assignment statements can only be used on type "reg" and need to be of the "non-blocking" type: <=
//always @(y) begin
//bird_y <= y;
//end


always @(posedge dclk or posedge clr)
begin

    if (!pause) begin

	    if (!gamestate && flap) gamestate = 1;
    
	    counter <= counter+1;
    
	    if (gamestate && counter % 200000 == 0) begin
		    if (flap) velocity <= 10;
		    else if (velocity < 20) velocity <= velocity + 1;
		
		    if (bird_y + velocity > 5 && bird_y + velocity < 455) bird_y <= bird_y + velocity;
	    end
    end
    
    
	// reset condition
	if (clr == 1)
	begin
		hc <= 0;
		vc <= 0;
		bird_y <= 10'd240;
		gamestate = 0;
		velocity <= -10;
	end
	else
	begin
		// keep counting until the end of the line
		if (hc < hpixels - 1)
			hc <= hc + 1;
		else
		// When we hit the end of the line, reset the horizontal
		// counter and increment the vertical counter.
		// If vertical counter is at the end of the frame, then
		// reset that one too.
		begin
			hc <= 0;
			if (vc < vlines - 1)
				vc <= vc + 1;
			else
				vc <= 0;
		end
		
	end
end

// generate sync pulses (active low)
// ----------------
// "assign" statements are a quick way to
// give values to variables of type: wire
assign hsync = (hc < hpulse) ? 0:1;
assign vsync = (vc < vpulse) ? 0:1;

// display 100% saturation colorbars
// ------------------------
// Combinational "always block", which is a block that is
// triggered when anything in the "sensitivity list" changes.
// The asterisk implies that everything that is capable of triggering the block
// is automatically included in the sensitivty list.  In this case, it would be
// equivalent to the following: always @(hc, vc)
// Assignment statements can only be used on type "reg" and should be of the "blocking" type: =
always @(*)
begin
	// first check if we're within vertical active video range
	if (vc >= vbp && vc < vfp)
	begin
		// now display different colors every 80 pixels
		// while we're within the active horizontal range
		// -----------------
		// display blue
		if (hc >= hbp && hc < (hbp+bird_x))
		begin
			red = 3'b000;
			green = 3'b101;
			blue = 3'b111;
		end
		// display yellow bar
		else if (hc >= (hbp+bird_x) && hc < (hbp+bird_x+20))
		begin
			if (vc >= (vbp+bird_y) && vc < (vbp+bird_y+20))
				begin
				// black part of the eyeball
				if (hc >= (hbp+bird_x+17) && hc < (hbp+bird_x+19) && vc >= (vbp+bird_y+13) && vc < (vbp+bird_y+15)) begin
					red = 0;
					green = 0;
					blue = 0;
				end
				// white part of the eyeball
				else if (hc >= (hbp+bird_x+15) && hc < (hbp+bird_x+20) && vc >= (vbp+bird_y+11) && vc < (vbp+bird_y+17)) begin
					red = 3'b111;
					green = 3'b111;
					blue = 3'b111;
				end 
				//rest of the bird
				else begin
					red = 3'b111;
					green = 3'b111;
					blue = 3'b000;
                  	end 
			// rest of the column	
			else begin
                      		red = 3'b000;
                      		green = 3'b100;
                      		blue = 3'b111;
                  	end
		end
		// display blue
		else if (hc >= (hbp+bird_x+20) && hc < (hfp))
		begin
			red = 3'b000;
			green = 3'b101;
			blue = 3'b111;
		end
		// we're outside active horizontal range so display black
		else
		begin
			red = 0;
			green = 0;
			blue = 0;
		end
	end
	// we're outside active vertical range so display black
	else
	begin
		red = 0;
		green = 0;
		blue = 0;
	end
	end
endmodule
